`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2020/11/10 15:47:21
// Design Name: 
// Module Name: controller
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//To generate instructions, shall be reformed to a decoder later
module controller(
    input clk,
    input rst,
    output wire[11:0]instruction,
    output reg[3:0][7:0]data//remember to remove this
    );
    reg psum_rst;
    assign instruction[0] = psum_rst;
    reg[3:0] bpug_sel;
    assign instruction[4:1] = bpug_sel;
    reg psum_add;
    assign instruction[5] = psum_add;
    reg img_data_sel;
    assign instruction[6] = img_data_sel;
    wire[1:0]en;
    assign instruction[8:7] = en;
    //reg[3:0]bpug_1sel;
    //assign instruction[11:8]=bpug_1sel;
    reg bpug_psum_add;
    assign instruction[9]=bpug_psum_add;
    reg cal_bin_wr;
    assign instruction[10]=cal_bin_wr;
    reg bias_wr;
    assign instruction[11] = bias_wr;
    
    reg[3:0] img_col;//col of image
    reg img_row;
    
    reg [7:0] cnt;
    reg if_cal;//if_cal==0, prepare data; if_cal==1, calculate
    reg [1:0]data_sel;//=2, image; =1, bias; =0, wgt
    wire [5:0]tesssst = {bpug_sel,2'b10};
    
    always@(posedge clk) begin
        if(rst) begin
            cnt <= 0;
            bpug_sel <= 0;
            if_cal<=0;
            data_sel <= 0;
            img_col <=0;
            img_row <=0;
        end
        else if(data_sel==2'b00)begin//read weight process
            if(cnt<6'b111011) cnt <= cnt+1'b1;
            else if(cnt==6'b111011) begin
                cnt <= 0;
                if(bpug_sel<2'b11) bpug_sel <= bpug_sel +1'b1;
                else if(bpug_sel == 2'b11) begin
                    bpug_sel <= 0;
                    data_sel <= 2'b01;//time to write bias data
                end
            end
        end
        
        else if(data_sel==2'b01)begin//writing bias
            if(cnt<4'b1101)begin
                cnt <= cnt+1'b1;
            end
            else if(cnt==4'b1101)begin
                cnt<=0;
                data_sel <=2'b10;
            end
        end
        
        //write image & calculation
        else if(data_sel==2'b10)begin
            if(cnt<60) begin
                cnt <= cnt+1'b1;
                if(img_col<6)begin
                    if(cnt==3)begin
                        cnt <= 0;
                        if(bpug_sel<2'b11) bpug_sel <= bpug_sel +1'b1;
                        else if(bpug_sel == 2'b11) begin
                            bpug_sel <= 0;
                            img_col <= img_col+1'b1;
                        end
                    end
                end
                else if(img_col>=6)begin
                    if(bpug_sel<2'b11) begin
                        if(cnt==3) begin
                            cnt <= 0;
                            bpug_sel <= bpug_sel +1'b1;
                        end
                    end
                end
            end
            else if(cnt==60) begin
                cnt <= 0;
                if(img_col<9) img_col <= img_col +1'b1;
                if(img_col==9) begin
                    img_col <= 0;
                    img_row <= ~img_row;
                end
            end
        end
    end
    
    reg wgt_en;
    assign en[0] = wgt_en;
    reg img_en;
    assign en[1] = img_en;

    wire[15:0][55:0][6:0] wgt;
    assign wgt = '{'{'{7'b0000011},'{7'b1011010},'{7'b0001000},'{7'b1011000},'{7'b1100100},'{7'b1000110},'{7'b1110000},'{7'b1000100},'{7'b1001000},'{7'b0000001},'{7'b1100010},'{7'b0111111},'{7'b0110110},'{7'b0011010},'{7'b0011011},'{7'b0001001},'{7'b0001000},'{7'b0011010},'{7'b0101110},'{7'b1011110},'{7'b1100110},'{7'b1110101},'{7'b0010111},'{7'b1110110},'{7'b1001100},'{7'b1001100},'{7'b0000001},'{7'b1110111},'{7'b0100010},'{7'b1110010},'{7'b1001000},'{7'b1110011},'{7'b0011001},'{7'b1100001},'{7'b1101001},'{7'b1100110},'{7'b0001101},'{7'b0001000},'{7'b0100110},'{7'b0111010},'{7'b0010011},'{7'b0000101},'{7'b1001101},'{7'b1111101},'{7'b0011110},'{7'b1011000},'{7'b1110010},'{7'b1011000},'{7'b0000000},'{7'b1110110},'{7'b0101000},'{7'b1100100},'{7'b1010010},'{7'b0011011},'{7'b1110110},'{7'b1110110}},'{'{7'b0001110},'{7'b0000110},'{7'b0000011},'{7'b0010000},'{7'b0000101},'{7'b1000011},'{7'b0011101},'{7'b1000110},'{7'b0000001},'{7'b1110100},'{7'b1011001},'{7'b1011010},'{7'b0101010},'{7'b0101110},'{7'b0001110},'{7'b0011101},'{7'b0011111},'{7'b0011111},'{7'b0101101},'{7'b0001011},'{7'b0001110},'{7'b1110101},'{7'b0101000},'{7'b0010000},'{7'b1101101},'{7'b1100001},'{7'b0110110},'{7'b0110001},'{7'b0011100},'{7'b0110010},'{7'b0000011},'{7'b0011100},'{7'b0010000},'{7'b1000101},'{7'b1001100},'{7'b1101010},'{7'b0111001},'{7'b0011010},'{7'b0111000},'{7'b0001100},'{7'b0011101},'{7'b1101000},'{7'b0000101},'{7'b0110101},'{7'b1110001},'{7'b0101110},'{7'b0000110},'{7'b0001110},'{7'b0101010},'{7'b1011011},'{7'b1100100},'{7'b0011001},'{7'b1100011},'{7'b0101010},'{7'b1001010},'{7'b1101100}},'{'{7'b0100000},'{7'b0101100},'{7'b1001001},'{7'b0000100},'{7'b0100010},'{7'b0001011},'{7'b0000111},'{7'b1111100},'{7'b1100000},'{7'b1110111},'{7'b0101111},'{7'b1010110},'{7'b1010011},'{7'b0011000},'{7'b0110010},'{7'b1111011},'{7'b1101000},'{7'b0100000},'{7'b1100001},'{7'b0001100},'{7'b1011100},'{7'b1101011},'{7'b0010101},'{7'b1010000},'{7'b0110000},'{7'b0000100},'{7'b1000000},'{7'b1011001},'{7'b1101011},'{7'b1011001},'{7'b0010010},'{7'b0010011},'{7'b0101010},'{7'b0000110},'{7'b1011001},'{7'b1000101},'{7'b0011011},'{7'b0011001},'{7'b0110110},'{7'b1110100},'{7'b0111010},'{7'b1111101},'{7'b0110000},'{7'b1001011},'{7'b1110011},'{7'b1100100},'{7'b0111010},'{7'b0100010},'{7'b1000000},'{7'b1011010},'{7'b0011011},'{7'b1101110},'{7'b1011101},'{7'b1010100},'{7'b1111100},'{7'b1011000}},'{'{7'b0100110},'{7'b0100110},'{7'b1001001},'{7'b0110011},'{7'b0110000},'{7'b1000111},'{7'b0000101},'{7'b1100101},'{7'b0001011},'{7'b1001110},'{7'b1101110},'{7'b0010110},'{7'b0101110},'{7'b1001111},'{7'b0001101},'{7'b1010111},'{7'b1010110},'{7'b0110111},'{7'b1011111},'{7'b1110010},'{7'b1001111},'{7'b1101100},'{7'b1000010},'{7'b0111000},'{7'b1010100},'{7'b1101011},'{7'b1100100},'{7'b1101110},'{7'b1011000},'{7'b1000000},'{7'b0101101},'{7'b1101100},'{7'b0011100},'{7'b0001100},'{7'b0000100},'{7'b0100001},'{7'b1100100},'{7'b0011001},'{7'b1101111},'{7'b1110111},'{7'b1001000},'{7'b1011101},'{7'b0000001},'{7'b0000101},'{7'b1110101},'{7'b0010101},'{7'b0010101},'{7'b0100110},'{7'b1110011},'{7'b0000010},'{7'b1111011},'{7'b0111101},'{7'b0111101},'{7'b0000100},'{7'b0101101},'{7'b1001011}},'{'{7'b1111011},'{7'b0001111},'{7'b1011100},'{7'b0010010},'{7'b0001001},'{7'b1001111},'{7'b1001101},'{7'b1100100},'{7'b0101000},'{7'b1101011},'{7'b1010011},'{7'b1111010},'{7'b1011111},'{7'b0100101},'{7'b0010011},'{7'b1000101},'{7'b0111011},'{7'b0011100},'{7'b0110000},'{7'b1111000},'{7'b1101001},'{7'b1010100},'{7'b1011100},'{7'b1001110},'{7'b1111010},'{7'b0100000},'{7'b0100101},'{7'b1111100},'{7'b1111010},'{7'b1100011},'{7'b1110000},'{7'b1000110},'{7'b0100001},'{7'b0100001},'{7'b1111101},'{7'b0100011},'{7'b1111100},'{7'b1000110},'{7'b0011011},'{7'b0011111},'{7'b1010010},'{7'b1001101},'{7'b1010110},'{7'b1111010},'{7'b0001100},'{7'b1101000},'{7'b0111001},'{7'b1000101},'{7'b1111111},'{7'b1000110},'{7'b0111110},'{7'b1111011},'{7'b1011110},'{7'b0111111},'{7'b0101010},'{7'b1000111}},'{'{7'b1111000},'{7'b1000010},'{7'b1101110},'{7'b1001001},'{7'b0101111},'{7'b1100101},'{7'b1011101},'{7'b0101110},'{7'b0010000},'{7'b1110111},'{7'b0100011},'{7'b0011001},'{7'b1101110},'{7'b1001111},'{7'b1010001},'{7'b0101110},'{7'b1000100},'{7'b0110011},'{7'b1111110},'{7'b0011011},'{7'b1000101},'{7'b1000010},'{7'b0110010},'{7'b0000111},'{7'b1110011},'{7'b0010011},'{7'b1110100},'{7'b1100010},'{7'b1001000},'{7'b1001110},'{7'b1110011},'{7'b1001001},'{7'b0101001},'{7'b0110011},'{7'b1101101},'{7'b0011100},'{7'b1100001},'{7'b0101010},'{7'b1110111},'{7'b1110111},'{7'b0111001},'{7'b0110010},'{7'b0101100},'{7'b0001010},'{7'b1001110},'{7'b1011010},'{7'b0001010},'{7'b0110001},'{7'b1001011},'{7'b0011100},'{7'b1011110},'{7'b0011110},'{7'b1100000},'{7'b0001010},'{7'b1010010},'{7'b0001011}},'{'{7'b0011011},'{7'b1100110},'{7'b1000101},'{7'b0110001},'{7'b1101001},'{7'b0011000},'{7'b1101001},'{7'b1100101},'{7'b1010011},'{7'b0101011},'{7'b1001101},'{7'b1110010},'{7'b0011011},'{7'b0011100},'{7'b0110011},'{7'b0001000},'{7'b1010011},'{7'b0010110},'{7'b1000110},'{7'b1000011},'{7'b0101111},'{7'b1101101},'{7'b0110100},'{7'b1101100},'{7'b0011000},'{7'b1100111},'{7'b0010011},'{7'b1100000},'{7'b0011001},'{7'b0111111},'{7'b0010110},'{7'b1101110},'{7'b1010100},'{7'b1001101},'{7'b1000010},'{7'b0011011},'{7'b1111010},'{7'b0001001},'{7'b0110110},'{7'b1000001},'{7'b0100000},'{7'b1001001},'{7'b0001011},'{7'b1101000},'{7'b1110100},'{7'b0101101},'{7'b0111001},'{7'b1100000},'{7'b0110101},'{7'b0011110},'{7'b0100000},'{7'b0001111},'{7'b0010001},'{7'b1101110},'{7'b1000011},'{7'b1010111}},'{'{7'b0110010},'{7'b0011001},'{7'b1010101},'{7'b0000110},'{7'b0110101},'{7'b1111100},'{7'b1010100},'{7'b0001110},'{7'b1011111},'{7'b0110111},'{7'b1011100},'{7'b1010111},'{7'b0010011},'{7'b1111010},'{7'b1101000},'{7'b0101101},'{7'b0001111},'{7'b0011100},'{7'b0010100},'{7'b1110000},'{7'b1101000},'{7'b0100101},'{7'b1101001},'{7'b0111100},'{7'b1001110},'{7'b0101011},'{7'b0100000},'{7'b1111111},'{7'b1000100},'{7'b1011000},'{7'b0010010},'{7'b1100011},'{7'b0000000},'{7'b1100010},'{7'b1101100},'{7'b0011100},'{7'b1000110},'{7'b1101101},'{7'b0111011},'{7'b0010110},'{7'b0001111},'{7'b1110000},'{7'b1100100},'{7'b1000100},'{7'b0111011},'{7'b0011100},'{7'b1010001},'{7'b1001010},'{7'b1011001},'{7'b1100000},'{7'b1101011},'{7'b0010011},'{7'b1010010},'{7'b1010110},'{7'b1010110},'{7'b1100001}},'{'{7'b1010011},'{7'b1101110},'{7'b0101110},'{7'b0110110},'{7'b0001100},'{7'b0100011},'{7'b1111111},'{7'b1001110},'{7'b0110001},'{7'b1101000},'{7'b0001011},'{7'b0111000},'{7'b0101011},'{7'b0000101},'{7'b0000010},'{7'b0110011},'{7'b1110111},'{7'b1111110},'{7'b1100010},'{7'b1000011},'{7'b0011100},'{7'b0001111},'{7'b1110101},'{7'b0110101},'{7'b1010010},'{7'b1100010},'{7'b0011011},'{7'b1010100},'{7'b0011101},'{7'b1101100},'{7'b1001000},'{7'b0000000},'{7'b0100111},'{7'b1000001},'{7'b1100101},'{7'b1110000},'{7'b1110011},'{7'b1101000},'{7'b1101111},'{7'b1111011},'{7'b1011000},'{7'b0100011},'{7'b0100000},'{7'b0110010},'{7'b1001111},'{7'b1101101},'{7'b1000001},'{7'b0111000},'{7'b1001001},'{7'b0011110},'{7'b1101111},'{7'b0000110},'{7'b1101001},'{7'b1100101},'{7'b0111001},'{7'b1011010}},'{'{7'b0100100},'{7'b0000100},'{7'b1100111},'{7'b0011111},'{7'b0101111},'{7'b0000110},'{7'b1111111},'{7'b1011111},'{7'b1001111},'{7'b0011100},'{7'b0101110},'{7'b1110111},'{7'b0001010},'{7'b0111100},'{7'b0011101},'{7'b0011111},'{7'b1100110},'{7'b1010011},'{7'b0100111},'{7'b0010110},'{7'b0111001},'{7'b0101011},'{7'b1110100},'{7'b0111110},'{7'b1000110},'{7'b0001010},'{7'b0111001},'{7'b1001111},'{7'b1101110},'{7'b0000100},'{7'b1110011},'{7'b1110010},'{7'b1000001},'{7'b0000001},'{7'b0100101},'{7'b0101100},'{7'b0100101},'{7'b0111000},'{7'b0011101},'{7'b0111110},'{7'b1010100},'{7'b0111110},'{7'b1000110},'{7'b1100010},'{7'b0101100},'{7'b1001111},'{7'b1000001},'{7'b1101101},'{7'b0001001},'{7'b0010110},'{7'b0100000},'{7'b0110001},'{7'b0100001},'{7'b1111111},'{7'b0111110},'{7'b0101111}},'{'{7'b0001101},'{7'b0101011},'{7'b1001101},'{7'b0110101},'{7'b0110111},'{7'b0000010},'{7'b1001010},'{7'b0001000},'{7'b1111110},'{7'b1001100},'{7'b0011000},'{7'b1101011},'{7'b0101000},'{7'b1110101},'{7'b1001100},'{7'b1011110},'{7'b0000010},'{7'b0111100},'{7'b0111101},'{7'b1101010},'{7'b1111010},'{7'b1001010},'{7'b0011101},'{7'b1011001},'{7'b1011111},'{7'b0011111},'{7'b1000101},'{7'b0111101},'{7'b1100110},'{7'b1001111},'{7'b0000111},'{7'b1101001},'{7'b1010101},'{7'b0110110},'{7'b0101101},'{7'b1011000},'{7'b0101010},'{7'b1101011},'{7'b1101100},'{7'b0011111},'{7'b1111100},'{7'b1111001},'{7'b1000001},'{7'b1110000},'{7'b1101010},'{7'b0110110},'{7'b0011100},'{7'b0001100},'{7'b0000010},'{7'b0000001},'{7'b0101101},'{7'b0111110},'{7'b0001110},'{7'b1001011},'{7'b1000010},'{7'b1010010}},'{'{7'b0010011},'{7'b1010001},'{7'b1000100},'{7'b0101011},'{7'b1001100},'{7'b0111100},'{7'b1000101},'{7'b0011111},'{7'b1110101},'{7'b0011001},'{7'b1111101},'{7'b0101100},'{7'b1010101},'{7'b0100010},'{7'b0101011},'{7'b1100001},'{7'b0011100},'{7'b1111001},'{7'b1001001},'{7'b1100101},'{7'b1100000},'{7'b0001001},'{7'b0101110},'{7'b0101110},'{7'b1001001},'{7'b1010010},'{7'b0001110},'{7'b1101101},'{7'b1100000},'{7'b0001110},'{7'b0011010},'{7'b0011111},'{7'b1110111},'{7'b1101000},'{7'b0101110},'{7'b1010001},'{7'b0011110},'{7'b1101010},'{7'b1111100},'{7'b1100100},'{7'b1000010},'{7'b0101000},'{7'b1100010},'{7'b0110010},'{7'b0100110},'{7'b1011000},'{7'b0100101},'{7'b0001010},'{7'b1001011},'{7'b0011000},'{7'b1000110},'{7'b0010011},'{7'b0101100},'{7'b1001111},'{7'b1011001},'{7'b0001101}},'{'{7'b0001100},'{7'b0100001},'{7'b1010101},'{7'b0100011},'{7'b0100111},'{7'b1011111},'{7'b1000100},'{7'b1000101},'{7'b0100011},'{7'b1001101},'{7'b1110100},'{7'b1010011},'{7'b1110110},'{7'b0010010},'{7'b1010111},'{7'b0011010},'{7'b0111111},'{7'b0100110},'{7'b0100111},'{7'b0110011},'{7'b1001010},'{7'b1101011},'{7'b0101110},'{7'b0000100},'{7'b0110100},'{7'b0010111},'{7'b0001100},'{7'b0010100},'{7'b1001111},'{7'b1100010},'{7'b1001001},'{7'b0010011},'{7'b0110111},'{7'b0100011},'{7'b1101101},'{7'b1111110},'{7'b1010000},'{7'b0011000},'{7'b0011000},'{7'b0110100},'{7'b1101111},'{7'b1000010},'{7'b0110111},'{7'b0101101},'{7'b0101101},'{7'b1011111},'{7'b1111110},'{7'b1110000},'{7'b1111000},'{7'b0111011},'{7'b0100011},'{7'b0111001},'{7'b1011111},'{7'b0000000},'{7'b0010100},'{7'b0111101}},'{'{7'b1000001},'{7'b1100010},'{7'b0010101},'{7'b1011011},'{7'b1010100},'{7'b1101000},'{7'b0101101},'{7'b1101011},'{7'b1010101},'{7'b0000101},'{7'b0001111},'{7'b0101100},'{7'b1101101},'{7'b0111100},'{7'b0111101},'{7'b0001011},'{7'b0111111},'{7'b1111100},'{7'b0011111},'{7'b1011000},'{7'b0011011},'{7'b0111111},'{7'b0101000},'{7'b0000000},'{7'b1011111},'{7'b1100101},'{7'b0100100},'{7'b1101010},'{7'b0110110},'{7'b1110101},'{7'b0000011},'{7'b1010101},'{7'b0101001},'{7'b1110000},'{7'b0010011},'{7'b0110010},'{7'b0001011},'{7'b1110101},'{7'b0000100},'{7'b1101100},'{7'b0110111},'{7'b0010111},'{7'b1001000},'{7'b0111110},'{7'b0111101},'{7'b0101101},'{7'b1111101},'{7'b1101000},'{7'b0100000},'{7'b0101000},'{7'b1010100},'{7'b0101001},'{7'b1000011},'{7'b0100001},'{7'b0111010},'{7'b1100100}},'{'{7'b1001111},'{7'b0000110},'{7'b1000100},'{7'b1101111},'{7'b1101000},'{7'b1111000},'{7'b1110000},'{7'b0011100},'{7'b0010010},'{7'b0010011},'{7'b0100100},'{7'b0011111},'{7'b1001110},'{7'b0101111},'{7'b1111110},'{7'b1100001},'{7'b1100000},'{7'b0100010},'{7'b1001110},'{7'b0100111},'{7'b0100100},'{7'b1010110},'{7'b1110010},'{7'b0100100},'{7'b1010000},'{7'b0111000},'{7'b1001111},'{7'b0101001},'{7'b1010001},'{7'b1011111},'{7'b1100011},'{7'b0111101},'{7'b1100000},'{7'b0101100},'{7'b1110001},'{7'b1111001},'{7'b0010001},'{7'b0011010},'{7'b1111011},'{7'b1110111},'{7'b1000001},'{7'b1100101},'{7'b0110100},'{7'b0000000},'{7'b0110000},'{7'b0100000},'{7'b0001011},'{7'b0100011},'{7'b1010010},'{7'b1100110},'{7'b1100101},'{7'b1010010},'{7'b1100100},'{7'b0111100},'{7'b0110001},'{7'b1111110}},'{'{7'b0000000},'{7'b0011011},'{7'b1011001},'{7'b0111000},'{7'b1101001},'{7'b0010000},'{7'b1101100},'{7'b0000000},'{7'b1111010},'{7'b1011000},'{7'b0010000},'{7'b0110010},'{7'b0000110},'{7'b1011011},'{7'b1000101},'{7'b0000110},'{7'b1100001},'{7'b1100001},'{7'b1101001},'{7'b0101101},'{7'b1110110},'{7'b0000111},'{7'b1110001},'{7'b1000100},'{7'b0010001},'{7'b0110010},'{7'b0010011},'{7'b1011000},'{7'b0001110},'{7'b1010011},'{7'b0100011},'{7'b0001110},'{7'b1101110},'{7'b1001011},'{7'b1110100},'{7'b1100011},'{7'b0111001},'{7'b0010001},'{7'b1101101},'{7'b0001110},'{7'b1001110},'{7'b0000110},'{7'b1001010},'{7'b1010101},'{7'b0001110},'{7'b0001011},'{7'b1000001},'{7'b0000010},'{7'b0100000},'{7'b0001100},'{7'b1111001},'{7'b0000000},'{7'b0110001},'{7'b1100000},'{7'b0001111},'{7'b0110000}}};

    always@(posedge clk) begin
        if(rst) begin
            wgt_en<=0;
        end
        else begin
            if(data_sel==2'b00) begin
                if(cnt<=6'b110111) begin
                    data[0]<=wgt[{bpug_sel,2'b00}][cnt];
                    data[1]<=wgt[{bpug_sel,2'b01}][cnt];
                    data[2]<=wgt[{bpug_sel,2'b10}][cnt];
                    data[3]<=wgt[{bpug_sel,2'b11}][cnt];
                    wgt_en <=1;
                end
                else if(cnt == 6'b111000)begin
                    wgt_en <= 0;
                end
            end
        end
    end
    
    wire[7:0][7:0]bias;
    assign bias = '{'{8'b11001000},'{8'b00001010},'{8'b01000110},'{8'b11010010},'{8'b10100100},'{8'b11001110},'{8'b01000000},'{8'b00101010}};
    always@(posedge clk)begin
        if(rst) begin
            bias_wr <= 0;
        end
        else if(data_sel==2'b01)begin
            if(cnt<=1'b1)begin
                data<={bias[{cnt,2'b00}],bias[{cnt,2'b01}],bias[{cnt,2'b10}],bias[{cnt,2'b11}]};
                bias_wr<=1;
            end
            else if(cnt==2'b10)begin
                bias_wr<=0;
            end
        end
    end
    wire[15:0][9:0][9:0] img_reg;
    assign img_reg ='{'{'{10'b0101100100},'{10'b1001100100},'{10'b1111100010},'{10'b1001110101},'{10'b1001100101},'{10'b0010110101},'{10'b1011011101},'{10'b1001111110},'{10'b0100001101},'{10'b0000000110}},
                    '{'{10'b0001010000},'{10'b0001010011},'{10'b1111000000},'{10'b1110100001},'{10'b0111101100},'{10'b0110110010},'{10'b0111000011},'{10'b1100010000},'{10'b1000001110},'{10'b0000000011}},
                    '{'{10'b1111001111},'{10'b1001111110},'{10'b0001101100},'{10'b0011000111},'{10'b0011010000},'{10'b1111111100},'{10'b1100100100},'{10'b0000001101},'{10'b0001001110},'{10'b0010100000}},
                    '{'{10'b0110011000},'{10'b0001101100},'{10'b0011010000},'{10'b0000011101},'{10'b0101000010},'{10'b1101100011},'{10'b0001100011},'{10'b1110011111},'{10'b0111001110},'{10'b1011001111}},
                    '{'{10'b0001101100},'{10'b0111001000},'{10'b0101000001},'{10'b1011111101},'{10'b1011101000},'{10'b1111111110},'{10'b0001010011},'{10'b0000010100},'{10'b0000000001},'{10'b1100001101}},
                    '{'{10'b1110101110},'{10'b0001011001},'{10'b1000001101},'{10'b1100110101},'{10'b1100010100},'{10'b1100110000},'{10'b1101111101},'{10'b0100000001},'{10'b1100010001},'{10'b0110000101}},
                    '{'{10'b1100100101},'{10'b0101010011},'{10'b1111000111},'{10'b1110111101},'{10'b1000111011},'{10'b0110001001},'{10'b0001111001},'{10'b0010001010},'{10'b0111110011},'{10'b1001011101}},
                    '{'{10'b0010000111},'{10'b0011001100},'{10'b0010111010},'{10'b1001011000},'{10'b0011000100},'{10'b1111001011},'{10'b1000100000},'{10'b0001001111},'{10'b0001011100},'{10'b1110110010}},
                    '{'{10'b0100011101},'{10'b1000010111},'{10'b0101100001},'{10'b0010101111},'{10'b0110001010},'{10'b1100000010},'{10'b1011001111},'{10'b1100001100},'{10'b1100001110},'{10'b1100010011}},
                    '{'{10'b0100001000},'{10'b0010001010},'{10'b0001111110},'{10'b0010100001},'{10'b1000111100},'{10'b1100110010},'{10'b0111100000},'{10'b1111001100},'{10'b1001111011},'{10'b0001111001}},
                    '{'{10'b1001000010},'{10'b0100010011},'{10'b1101010010},'{10'b0010110101},'{10'b1111000100},'{10'b0100100101},'{10'b0001110010},'{10'b1001101110},'{10'b0111011111},'{10'b1101011010}},
                    '{'{10'b0110010111},'{10'b0101110100},'{10'b1100000111},'{10'b1101101100},'{10'b1011001101},'{10'b1101000110},'{10'b0110101111},'{10'b1000011100},'{10'b0111001110},'{10'b0110110000}},
                    '{'{10'b0001010011},'{10'b0101111001},'{10'b1110101011},'{10'b0101001011},'{10'b1110010100},'{10'b0101000110},'{10'b0001100101},'{10'b0011110000},'{10'b1010011111},'{10'b1011000000}},
                    '{'{10'b1111011011},'{10'b1011100011},'{10'b0101001000},'{10'b0100101101},'{10'b0010000011},'{10'b0100010110},'{10'b1010111000},'{10'b0000100000},'{10'b1100000010},'{10'b0000010111}},
                    '{'{10'b0101000000},'{10'b0110000011},'{10'b0011010111},'{10'b0010000111},'{10'b0001000111},'{10'b1110110111},'{10'b1000110010},'{10'b1110000100},'{10'b1011000001},'{10'b0100010110}},
                    '{'{10'b1100011101},'{10'b0011011001},'{10'b0010101011},'{10'b0100100010},'{10'b0011010100},'{10'b0011101100},'{10'b1000001000},'{10'b0001100010},'{10'b1101101100},'{10'b0011101011}}};
    
    wire [3:0][7:0]fxx_k;
    wire[3:0][5:0] bpug_sel_extend = {{bpug_sel,2'b11},{bpug_sel,2'b10},{bpug_sel,2'b01},{bpug_sel,2'b00}}; 
    assign fxx_k[0] = img_reg[bpug_sel_extend[0]][img_col]>>(2*img_row);//{img_reg[bpug_sel_extend[3]][img_col]>>(2*img_row),img_reg[bpug_sel_extend[2]][img_col]>>(2*img_row),img_reg[bpug_sel_extend[1]][img_col]>>(2*img_row),};
    assign fxx_k[1] = img_reg[bpug_sel_extend[1]][img_col]>>(2*img_row);
    assign fxx_k[2] = img_reg[bpug_sel_extend[2]][img_col]>>(2*img_row);
    assign fxx_k[3] = img_reg[bpug_sel_extend[3]][img_col]>>(2*img_row);
    always@(posedge clk) begin
        if(rst) begin
            img_en<=0;
        end
        else if(data_sel==2'b10)begin
            if(cnt==1) begin
                data<=fxx_k;
                img_en <=1;
            end
            else if(cnt == 2)begin
                img_en <= 0;
            end
        end
    end
    
    always@(posedge clk) begin
        if(rst) begin
            bpug_sel <= 0;
            psum_rst <= 0;
            psum_add <= 0;
            bpug_psum_add<=0;
            img_data_sel <= 0;
            cal_bin_wr<= 0;
        end
        else if(data_sel==2'b10) case(cnt)
            5: begin
                bpug_sel <= 0;//in this section bpug is used to select BPUE
                psum_rst <= 1;
                img_data_sel <= 0;
            end
            6:begin
                psum_rst <= 0;
            end
            7:begin
                psum_add <=1;
                bpug_sel <= 1;
            end
            8:begin
                bpug_sel <= 2;
            end
            9:begin
                bpug_sel <= 3; 
            end
            10:begin
                bpug_sel <= 4;
            end
            11:begin
                bpug_sel <= 5;
            end
            12:begin
                bpug_sel <= 6;
            end
            14:begin
                psum_add<=0;
                bpug_sel <= 0;
            end
            
            15:begin
                bpug_psum_add <= 1;
                bpug_sel<=0;//in this section bpug is used to select BPUG
            end
            16:begin
                bpug_sel<=1;
            end
            17:begin
                bpug_sel<=2;
            end
            18:begin
                bpug_sel<=3;
            end
            19:begin
                bpug_sel<=4;
            end
            20:begin
                bpug_sel<=5;
            end
            21:begin
                bpug_sel<=6;
            end
            22:begin
                bpug_sel<=7;
            end
            23:begin
                bpug_sel<=8;
            end
            24:begin
                bpug_sel<=9;
            end
            25:begin
                bpug_sel<=10;
            end
            26:begin
                bpug_sel<=11;
            end
            27:begin
                bpug_sel<=12;
            end
            28:begin
                bpug_sel<=13;
            end
            29:begin
                bpug_sel<=14;
            end
            30:begin
                bpug_sel <= 15;
            end
            31:begin
                bpug_psum_add <= 0;
                bpug_sel <= 0;
                cal_bin_wr<=1;
            end
            32:begin
                cal_bin_wr<=0;
                psum_rst <= 1;
                img_data_sel <= 1;
            end
            33:begin
                psum_rst <= 0;
            end
            34:begin
                psum_add <=1;
                bpug_sel <= 1;//again BPUE
            end
            35:begin
                bpug_sel <= 2;
            end
            36:begin
                bpug_sel <= 3; 
            end
            37:begin
                bpug_sel <= 4;
            end
            38:begin
                bpug_sel <= 5;
            end
            39:begin
                bpug_sel <= 6;
            end
            41:begin
                psum_add<=0;
                bpug_sel <= 0;
            end

            42:begin
                bpug_psum_add <= 1;
                bpug_sel<=0;
            end
            43:begin
                bpug_sel<=1;
            end
            44:begin
                bpug_sel<=2;
            end
            45:begin
                bpug_sel<=3;
            end
            46:begin
                bpug_sel<=4;
            end
            47:begin
                bpug_sel<=5;
            end
            48:begin
                bpug_sel<=6;
            end
            49:begin
                bpug_sel<=7;
            end
            50:begin
                bpug_sel<=8;
            end
            51:begin
                bpug_sel<=9;
            end
            52:begin
                bpug_sel<=10;
            end
            53:begin
                bpug_sel<=11;
            end
            54:begin
                bpug_sel<=12;
            end
            55:begin
                bpug_sel<=13;
            end
            56:begin
                bpug_sel<=14;
            end
            57:begin
                bpug_sel <= 15;
            end
            58:begin
                bpug_psum_add <= 0;
                bpug_sel <= 0;
                cal_bin_wr<=1;
            end
            59:begin
                cal_bin_wr<=0;
            end
        endcase
    end
endmodule
